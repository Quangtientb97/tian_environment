// --------------------------------------------
// File Name   : reg_pkg.sv
// Description :
// Developers  :
// Created     :
// Generator   : csv_regdef
// --------------------------------------------

`ifndef SUV_REG_PKG
`define SUV_REG_PKG

//--------------------------------------------------------
//  BE CAREFUL CHANGING FOLLOWING IMPORT ORDER! 
//--------------------------------------------------------
//--------------------------------------------------------
//  Import UVM library macros.
//--------------------------------------------------------
`include "uvm_macros.svh"

//--------------------------------------------------------
//  Include macros. 
//--------------------------------------------------------
`include "reg_def_defines.sv"

package reg_pkg;
	//--------------------------------------------------------
	//  Import UVM library 
	//--------------------------------------------------------
	import uvm_pkg::*;

	//--------------------------------------------------------
	//  Include register of each IP 
	//--------------------------------------------------------
	__INCLUDE_REG_DEF_FILE__

	//--------------------------------------------------------
	//  Include register block of top 
	//--------------------------------------------------------
	`include "reg_blk.sv"

endpackage: reg_pkg

`endif //SUV_REG_PKG

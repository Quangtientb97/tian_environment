`define CLOCK_PERIOD 5
`define RESET_CYCLE 10

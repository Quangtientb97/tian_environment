`ifndef ADDR_WIDTH
	`define ADDR_WIDTH 8
`endif //ADDR_WIDTH

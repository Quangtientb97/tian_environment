// class seq0 extends seq_lib
// use `uvm_do and `uvm_do_with to excecute sequence
